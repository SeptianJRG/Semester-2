library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Post_Test is
	port(A,B : in STD_LOGIC_VECTOR(1 downto 0);
		x,y,z : out STD_LOGIC);
	
end Post_Test;

architecture Behavioral of Post_Test is

begin
	

end Behavioral;

