library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity fire_alarm is
	fire: in std_logic;
	fire_sensor:
	arm_disarm_btn
	
end fire_alarm;

architecture Behavioral of fire_alarm is

begin


end Behavioral;

